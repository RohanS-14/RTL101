//clock buffer
module clkbuff(input iclk,output oclk);

buf b1(oclk,iclk);

endmodule
