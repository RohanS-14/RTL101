module couter_tb1();
reg clk,rst,load;
wire [0:3] q;
reg [0:3] dn;